import os;import net.http;const list_url = "https://raw.githubusercontent.com/watakak/VLib/refs/heads/main/list.txt";const modules_dir=os.home_dir()+"\\.vmodules";fn fetch_module_list()map[string]string{response:=http.get(list_url)or{eprintln("Failed to fetch the module list: $err");return{}};mut modules:=map[string]string{};for line in response.body.split("\n"){if line.trim_space().len==0||line.starts_with("#"){continue};parts:=line.split(" ");if parts.len==2{modules[parts[0]]=parts[1].trim_right("/")}};return modules};fn install_module(name string,url string)!{if!os.exists(modules_dir){os.mkdir(modules_dir)!};dest_dir:=os.join_path(modules_dir,name);if os.exists(dest_dir){println("Module '$name' is already installed.");return};println("Downloading module '$name' from $url");zip_path:=dest_dir+".zip";println(".zip file path: $zip_path");http.download_file(url+"/archive/refs/heads/main.zip",zip_path)!;if!os.exists(zip_path){return error("Download completed but zip file not found: $zip_path")};zip_size:=os.file_size(zip_path);println("Downloaded .zip file size: $zip_size bytes");temp_dir:=os.join_path(modules_dir,"temp_extraction");os.mkdir(temp_dir)!;extraction_result:=os.execute("powershell -Command \"Expand-Archive -Path '${zip_path}' -DestinationPath '${temp_dir}'\"");if extraction_result.exit_code!=0{os.rmdir_all(temp_dir)!;return error("Failed to extract module archive: ${extraction_result.output}")};entries:=os.ls(temp_dir)or{os.rmdir_all(temp_dir)!;return error("Failed to list contents of the temporary extraction directory: $err")};if entries.len==0{os.rmdir_all(temp_dir)!;return error("No files or directories found in the extracted archive.")};original_dir:=os.join_path(temp_dir,entries[0]);if!os.is_dir(original_dir){os.rmdir_all(temp_dir)!;return error("Expected a directory but found something else: ${original_dir}")};os.mv(original_dir,dest_dir)!;os.rmdir_all(temp_dir)!;os.rm(zip_path)!;println("Module '$name' has been successfully installed.")};fn uninstall_module(name string)!{dest_dir:=os.join_path(modules_dir,name);if!os.exists(dest_dir){println("Module '$name' is not installed.");return};println("Removing module directory: $dest_dir");os.rmdir_all(dest_dir)!;println("Module '$name' has been successfully uninstalled.")};fn main(){if os.args.len<3{println("Usage: vlib <command> <module_name>");return};command:=os.args[1];module_name:=os.args[2];modules:=fetch_module_list();match command{"install"{if module_name!in modules{println("Module '$module_name' not found in the list.");return};install_module(module_name,modules[module_name])or{eprintln("Error: $err")}}"uninstall"{uninstall_module(module_name)or{eprintln("Error: $err")}}else{println("Unknown command: $command");println("Usage: vlib <install|uninstall> <module_name>")}}}
